
/* Memoria ROM 8 Bits
INPUTS:
address: Posición de memoria van de 4 en 4
OUTPUTS
data: Valor almacenado de 8 bits
*/
module ROM8(
	input logic[10:0] address, 
	output logic[7:0] data
	);
	always @*
		case(address)
			11'h000: data = 8'b00000001; //
			11'h001: data = 8'b00000000; //
			11'h002: data = 8'b00000000; //
			11'h003: data = 8'b00000000; //
			11'h004: data = 8'b00000000; //
			11'h005: data = 8'b00000000; //
			11'h006: data = 8'b00000000; //
			11'h007: data = 8'b00000000; //
			11'h008: data = 8'b00000000; //
			11'h009: data = 8'b00000000; //
			11'h00a: data = 8'b00000000; //
			11'h00b: data = 8'b00000000; //
			11'h00c: data = 8'b00000000; //
			11'h00d: data = 8'b00000000; //
			11'h00f: data = 8'b00000000; //
		
			11'h010: data = 8'b00000001; //
			11'h011: data = 8'b00000000; //
			11'h012: data = 8'b00000000; //
			11'h013: data = 8'b00000000; //
			11'h014: data = 8'b00000000; //
			11'h015: data = 8'b00000000; //
			11'h016: data = 8'b00000000; //
			11'h017: data = 8'b00000000; //
			11'h018: data = 8'b00000000; //
			11'h019: data = 8'b00000000; //
			11'h01a: data = 8'b00000000; //
			11'h01b: data = 8'b00000000; //
			11'h01c: data = 8'b00000000; //
			11'h01d: data = 8'b00000000; //
			11'h01f: data = 8'b00000000; //
			
			11'h020: data = 8'b00000001; //
			11'h021: data = 8'b00000000; //
			11'h022: data = 8'b00000000; //
			11'h023: data = 8'b00000000; //
			11'h024: data = 8'b00000000; //
			11'h025: data = 8'b00000000; //
			11'h026: data = 8'b00000000; //
			11'h027: data = 8'b00000000; //
			11'h028: data = 8'b00000000; //
			11'h029: data = 8'b00000000; //
			11'h02a: data = 8'b00000000; //
			11'h02b: data = 8'b00000000; //
			11'h02c: data = 8'b00000000; //
			11'h02d: data = 8'b00000000; //
			11'h02f: data = 8'b00000000; //
			
			11'h030: data = 8'b00000001; //
			11'h031: data = 8'b00000000; //
			11'h032: data = 8'b00000000; //
			11'h033: data = 8'b00000000; //
			11'h034: data = 8'b00000000; //
			11'h035: data = 8'b00000000; //
			11'h036: data = 8'b00000000; //
			11'h037: data = 8'b00000000; //
			11'h038: data = 8'b00000000; //
			11'h039: data = 8'b00000000; //
			11'h03a: data = 8'b00000000; //
			11'h03b: data = 8'b00000000; //
			11'h03c: data = 8'b00000000; //
			11'h03d: data = 8'b00000000; //
			11'h03f: data = 8'b00000000; //
			
			
			default: data = 8'b00000000;
			
			
		endcase 
	
		
	
endmodule 