/* 
	Memoria de datos.
	Contiene las palabras descifradas. Los últimos 8 bits (LSB) Contienen el valor de la palbra.
*/

module dataMemory(input logic clk,
					input logic we, 	//Señal de Write Enable (permitir escritura)
					input logic[7:0] address, //posición de memoria -> 0 - 255 -> 2^8
					input logic [31:0] wdata, //Write data value -> Write value port
					output logic [31:0] rdata);//Read data value -> read value port 
	
	logic [7:0] RAM[255:0]; //255 celdas de 8-bit cada uno de ellas. Cada celda se accede de la forma: RAM[<numeroDelaCelda>]

	
	
	//Para la ESCRITURA en la memoria unicamente cuando se de el posedge del CLK y el enable este en 1.
	always_ff @(posedge clk)
		if (we) {RAM[address],RAM[address+1], RAM[address+2], RAM[address+3] } <= wdata;
		
	//Para la LECTURA del contenido en la RAM. 
	assign rdata = (we == 1'b0) ? {RAM[address],RAM[address+1], RAM[address+2], RAM[address+3]}  : 32'b0; //Si no se está haciendo una potencial escritura(Write Enable = 1), tomar la dirección a la que se apunta en address.
	
endmodule